interface rstn_if (input logic clk);
 logic rstn;
endinterface : rstn_if