interface clk_if();

    logic clk;

endinterface : clk_if